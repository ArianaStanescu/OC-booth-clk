module booth(
  input clk, bgn, rst
);
