module xor_m_3( 
  input wire m, c3,
  output wire out);
  
  
  assign out = m ^ c3;

endmodule

