library verilog;
use verilog.vl_types.all;
entity adder_xor_tb is
end adder_xor_tb;
