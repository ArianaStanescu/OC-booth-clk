library verilog;
use verilog.vl_types.all;
entity xor_m_c3 is
    port(
        m               : in     vl_logic;
        c3              : in     vl_logic;
        \out\           : out    vl_logic
    );
end xor_m_c3;
