library verilog;
use verilog.vl_types.all;
entity xor_gate_tb is
end xor_gate_tb;
